module tb_linx_cpu_pyc;
  logic clk;
  logic rst;

  logic [63:0] boot_pc = 64'h0000_0000_0001_0000;
  logic [63:0] boot_sp = 64'h0000_0000_0002_0000;

  logic halted;
  logic [63:0] pc;
  logic [2:0] stage;
  logic [63:0] cycles;
  logic [63:0] a0;
  logic [63:0] a1;
  logic [63:0] ra;
  logic [63:0] sp;
  logic [1:0] br_kind;
  logic [63:0] if_window;
  logic [5:0] wb_op;
  logic [5:0] wb_regdst;
  logic [63:0] wb_value;
  logic commit_cond;
  logic [63:0] commit_tgt;

  // Generated by pyc-compile: module linx_cpu_pyc
  linx_cpu_pyc dut (
      .clk(clk),
      .rst(rst),
      .boot_pc(boot_pc),
      .boot_sp(boot_sp),
      .halted(halted),
      .pc(pc),
      .stage(stage),
      .cycles(cycles),
      .a0(a0),
      .a1(a1),
      .ra(ra),
      .sp(sp),
      .br_kind(br_kind),
      .if_window(if_window),
      .wb_op(wb_op),
      .wb_regdst(wb_regdst),
      .wb_value(wb_value),
      .commit_cond(commit_cond),
      .commit_tgt(commit_tgt)
  );

  always #5 clk = ~clk;

  function automatic logic [31:0] mem_read32(input int unsigned addr);
    mem_read32 = {dut.mem.mem[addr + 3], dut.mem.mem[addr + 2], dut.mem.mem[addr + 1], dut.mem.mem[addr + 0]};
  endfunction

  string memh_path;
  int unsigned expected;
  string vcd_path;
  string log_path;
  int log_fd;
  bit log_cycles;
  int i;
  logic [31:0] got;

  initial begin
    clk = 1'b0;
    rst = 1'b1;
    if (!$value$plusargs("memh=%s", memh_path)) begin
      memh_path = "examples/linx_cpu/programs/test_or.memh";
    end
    if (!$value$plusargs("expected=%h", expected)) begin
      expected = 32'h0000_ff00;
    end

    // Tracing / logging (default: enabled; disable with +notrace / +nolog).
    vcd_path = "examples/generated/linx_cpu_pyc/tb_linx_cpu_pyc_sv.vcd";
    log_path = "examples/generated/linx_cpu_pyc/tb_linx_cpu_pyc_sv.log";
    void'($value$plusargs("vcd=%s", vcd_path));
    void'($value$plusargs("log=%s", log_path));
    log_cycles = $test$plusargs("logcycles");

    if (!$test$plusargs("notrace")) begin
      $display("tb_linx_cpu_pyc: dumping VCD to %s", vcd_path);
      $dumpfile(vcd_path);
      $dumpvars(0, tb_linx_cpu_pyc);
    end

    if (!$test$plusargs("nolog")) begin
      log_fd = $fopen(log_path, "w");
      $fdisplay(log_fd, "tb_linx_cpu_pyc(SV): memh=%s expected=0x%08x", memh_path, expected);
      $fdisplay(log_fd, "cycle,time,halted,stage,pc,cycles");
    end else begin
      log_fd = 0;
    end

    $display("tb_linx_cpu_pyc: memh=%s expected=0x%08x", memh_path, expected);

    $readmemh(memh_path, dut.mem.mem);

    repeat (5) @(posedge clk);
    rst = 1'b0;

    i = 0;
    while (i < 200000 && !halted) begin
      @(posedge clk);
      if (log_fd != 0 && log_cycles) begin
        $fdisplay(log_fd, "%0d,%0t,%0b,%0d,0x%016x,%0d", i, $time, halted, stage, pc, cycles);
      end
      i++;
    end

    if (!halted) begin
      $fatal(1, "FAIL: did not halt (pc=0x%016x cycles=%0d)", pc, cycles);
    end

    got = mem_read32(32'h0000_0100);
    if (got !== expected[31:0]) begin
      $fatal(1, "FAIL: mem[0x100]=0x%08x expected=0x%08x", got, expected[31:0]);
    end

    if (log_fd != 0) begin
      $fdisplay(log_fd, "PASS: mem[0x100]=0x%08x cycles=%0d pc=0x%016x", got, cycles, pc);
      $fclose(log_fd);
    end

    $display("PASS: mem[0x100]=0x%08x cycles=%0d", got, cycles);
    $finish;
  end

endmodule
